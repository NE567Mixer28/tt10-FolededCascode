** sch_path: /home/ttuser/tt10-FoldedCascode/xschem/untitled-4.sch
**.subckt untitled-4 VDD GND IN+
*.iopin VDD
*.iopin GND
*.ipin IN+
VbiasR1 IN+ net1 0 ac 1 0 sin(0 500u 50 0 0 0)
V2 net1 GND 0.9
V1 VDD GND 1.8
XM1 D IN+ VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XR5 GND Vc GND sky130_fd_pr__res_xhigh_po W=0.35 L=3.2 mult=1 m=1
XR2 Vc VDD GND sky130_fd_pr__res_xhigh_po W=0.35 L=5 mult=1 m=1
XR3 Vp VDD GND sky130_fd_pr__res_xhigh_po W=0.35 L=5 mult=1 m=1
XR4 GND Vp GND sky130_fd_pr__res_xhigh_po W=0.35 L=1.94 mult=1 m=1
**** begin user architecture code



.option reltol=1e-5
+  abstol=1e-14 savecurrents
.control
  save all
  op
  remzerovec
  write OTA_FoldedCascode_Noise.raw

  set appendwrite
  noise v(D) VbiasR1 dec 10 0.01 1e3
  remzerovec
  write OTA_FoldedCascode_Noise.raw

.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
