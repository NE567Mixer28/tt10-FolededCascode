** sch_path: /home/ttuser/tt10-FoldedCascode/xschem/retePmos.sch
**.subckt retePmos VDD GND
*.iopin VDD
*.iopin GND
XM7 G Vc2 D9 D9 sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 D9 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 D10 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 G Vc2 D10 D10 sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 VDD GND 1.8
V3 OUT GND 0.9
V5 Vc2 GND 0.45
I0 G GND 25u
I1 G GND 25u
**** begin user architecture code



* ngspice commands

.options savecurrents

.control
save all

save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm9.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]

   op
   remzerovec
   write retePmos.raw
   set appendwrite


.endc
.end




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
