** sch_path: /home/ttuser/tt10-FoldedCascode/xschem/ecg_pwl1_1.sch
**.subckt ecg_pwl1_1 VDD GND VDD VDD GND GND VDD GND VDD GND VDD GND VDD GND VDD GND VDD GND VDD GND VDD GND VDD GND VDD GND VDD
*+ GND VDD GND VDD GND VDD GND VDD GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin VDD
*.iopin GND
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
*.iopin VDD
*.iopin GND
V3 VDD GND 1.8
R1 net3 out1 250k m=1
R2 net4 out2 250k m=1
R6 net1 out_ref 250k m=1
R8 out net5 100k m=1
C1 out_ref net5 10u m=1
R5 net2 out 250k m=1
R4 out12 net2 10k m=1
R7 out22 net1 10k m=1
R9 net7 A 430k m=1
C2 ref net6 2.45n m=1
R10 net6 net7 430k m=1
C3 outPB net7 2.45n m=1
R11 ref net8 500k m=1
C5 net15 net9 4u m=1
C6 net9 net8 4u m=1
R13 outA net11 250k m=1
R14 net11 net12 10k m=1
R16 out_drl net13 220k m=1
R17 net13 net14 220 m=1
C4 net13 out_drl 100n m=1
C7 GND outPA 100n m=1
R18 outPA net10 100 m=1
R12 net9 net10 500k m=1
XR3 Vcm net3 GND sky130_fd_pr__res_high_po_0p35 L=0.4 mult=1 m=1
XR15 Vcm net4 GND sky130_fd_pr__res_high_po_0p35 L=0.4 mult=1 m=1
R19 net21 net20 302.1k m=1
R20 net17 net21 302.1k m=1
R21 net16 net18 151.05k m=1
C8 net21 net16 20n m=1
C9 net18 net20 10n m=1
C10 net17 net18 10n m=1
R22 net19 outN 100 m=1
R23 ref net19 100k m=1
x1 VDD GND out1 net3 IN1 OFC1_1
x2 VDD GND out2 net4 IN2 OFC1_1
x3 VDD GND out12 out12 out1 OFC1_1
x4 VDD GND out22 out22 out2 OFC1_1
x5 VDD GND out net2 net1 OFC1_1
x6 VDD GND out_ref net5 ref OFC1_1
x7 VDD GND net14 net14 Vcm OFC1_1
x8 VDD GND out_drl net13 ref OFC1_1
x9 VDD GND net12 net12 out OFC1_1
x10 VDD GND outA net11 ref OFC1_1
x11 VDD GND A A outA OFC1_1
x12 VDD GND outPB outPB net6 OFC1_1
x13 VDD GND net15 net15 outPB OFC1_1
x14 VDD GND net10 net10 net8 OFC1_1
x15 VDD GND net20 net20 outPA OFC1_1
x16 VDD GND outN outN net17 OFC1_1
x17 VDD GND net16 net16 net19 OFC1_1
**** begin user architecture code


** --- IMPOSTAZIONI DI SIMULAZIONE ---
.option reltol=1e-3 abstol=1e-12 method=gear

* --- DEFINIZIONE GENERATORI (Seguendo Immagine 2026-01-03 122450.png) ---

* V2: Generatore di Bias Principale (Offset 0.9V)
V2 v_offset GND 0.9

* VbiasR3: Generatore di MODO COMUNE (50Hz)
* Iniettato nel punto comune 'ref', sollevato dall'offset di 0.9V
VbiasR3 ref v_offset dc 0 sin(0 100m 50 0 0 0)

* VbiasR1: Braccio Positivo (ECG / 2)
* Collegato tra IN1 e ref. Fase 0.
VbiasR1 IN1 ref dc 0 pwl(
+ 0.00 0.00000 0.05 0.00000 0.08 0.00000 0.10 0.00005 0.12 0.000075
+ 0.15 0.00010 0.18 0.000075 0.22 0.00000 0.28 0.00000 0.29 -0.000025
+ 0.30 -0.00005 0.31 0.00035 0.32 0.00075 0.33 0.00035 0.34 -0.00010
+ 0.35 -0.00005 0.36 0.00000 0.40 0.00000 0.48 0.00000 0.52 0.00005
+ 0.56 0.000125 0.60 0.00015 0.64 0.000125 0.68 0.00005 0.75 0.00000
+ 1.00 0.00000 )

* VbiasR2: Braccio Negativo (ECG / 2 Invertito)
* Collegato tra IN2 e ref. I valori del PWL sono moltiplicati per -1.
VbiasR2 IN2 ref dc 0 pwl(
+ 0.00 0.00000 0.05 0.00000 0.08 0.00000 0.10 -0.00005 0.12 -0.000075
+ 0.15 -0.00010 0.18 -0.000075 0.22 0.00000 0.28 0.00000 0.29 0.000025
+ 0.30 0.00005 0.31 -0.00035 0.32 -0.00075 0.33 -0.00035 0.34 0.00010
+ 0.35 0.00005 0.36 0.00000 0.40 0.00000 0.48 0.00000 0.52 -0.00005
+ 0.56 -0.000125 0.60 -0.00015 0.64 -0.000125 0.68 -0.00005 0.75 0.00000
+ 1.00 0.00000 )

* --- CONTROLLO SIMULAZIONE ---
.control
    * Salvataggio segnali per analisi MATLAB
    save v(IN1) v(IN2) v(ref) v(outN)

    tran 10u 1.1s 0 1m

    * Plot per verifica differenziale
    * L'ECG utile è v(IN1)-v(IN2). Il rumore comune è v(ref)-0.9.
    plot v(IN1) v(IN2) title 'Ingressi OTA: IN1 e IN2 (Differenziali + Comune)'
    plot (v(IN1)-v(IN2)) title 'Segnale ECG Differenziale Puro'
    plot v(outN)
    * Esportazione dati (Tempo, IN1, IN2, Uscita)
    wrdata dati_ecg1.txt  v(outN)
.endc
.end




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  OFC1_1.sym # of pins=5
** sym_path: /home/ttuser/tt10-FoldedCascode/xschem/OFC1_1.sym
** sch_path: /home/ttuser/tt10-FoldedCascode/xschem/OFC1_1.sch
.subckt OFC1_1 VDD GND OUT IN- IN+
*.iopin VDD
*.iopin GND
*.ipin IN+
*.ipin IN-
*.opin OUT
XM11 S Vb VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=85 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM1 D1 IN+ S S sky130_fd_pr__pfet_01v8_lvt L=10 W=50 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 D2 IN- S S sky130_fd_pr__pfet_01v8_lvt L=10 W=50 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 OUT Vc1 D2 GND sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 D2 Vc GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 D1 Vc GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 G Vc1 D1 GND sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR2 Vb VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR3 GND Vb GND sky130_fd_pr__res_xhigh_po_0p35 L=13.2 mult=1 m=1
XR1 Vc VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR4 GND Vc GND sky130_fd_pr__res_xhigh_po_0p35 L=3.07 mult=1 m=1
XR5 Vc1 VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR6 GND Vc1 GND sky130_fd_pr__res_xhigh_po_0p35 L=13.2 mult=1 m=1
XR7 Vc2 VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR8 GND Vc2 GND sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XM7 G Vc2 D9 VDD sky130_fd_pr__pfet_01v8_lvt L=1.2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 D9 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1.2 W=5.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 D10 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1.2 W=5.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 OUT Vc2 D10 VDD sky130_fd_pr__pfet_01v8_lvt L=1.2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 OUT D1 sky130_fd_pr__cap_mim_m3_1 W=50 L=20 MF=1 m=1
.ends

.GLOBAL GND
.end
