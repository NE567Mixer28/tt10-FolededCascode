** sch_path: /home/ttuser/tt10-FoldedCascode/xschem/Pmos_noise.sch
**.subckt Pmos_noise VDD GND IN+
*.iopin VDD
*.iopin GND
*.ipin IN+
VbiasR1 IN+ net1 0 ac 1 0
V2 net1 GND 0.9
V1 VDD GND 1.8
C1 D GND 1p m=1
XM1 D IN+ S VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
V3 Vb GND 1.3
R1 D GND 70k m=1
XM3 S Vb VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=90 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM2 D1 IN- S VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
V4 IN- GND 0.9
R2 D1 GND 70k m=1
C2 D1 GND 1p m=1
**** begin user architecture code



.option reltol=1e-5
+  abstol=1e-14 savecurrents

.control

  save all
  save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]
  op
  remzerovec
  write Pmos_noise.raw

  set appendwrite
  noise v(D) VbiasR1 dec 10 0.1 100
  remzerovec
  write Pmos_noise.raw
  setplot noise1
  plot inoise_spectrum
  wrdata ~/Desktop/SIm/noise_W5.dat frequency inoise_spectrum

.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
